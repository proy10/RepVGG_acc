module mul #(
	parameter DW_IN = 8,
	parameter DW_OUT = 16
	)(
	input [DW_IN-1:0]	fmap,
	input [DW_IN-1:0]	wht,
	
	output [DW_OUT-1:0]	re
);
	
	

endmodule
