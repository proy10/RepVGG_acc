/*

*/

module pe(
	
);

endmodule
